library verilog;
use verilog.vl_types.all;
entity Coor_gen_tb is
end Coor_gen_tb;
